`include "logs.svh"








package packet_pkg;

    typedef bit [7:0] data_t[];



    class Packet;
        data_t      data;
        bit         err;
    
        function automatic int size();
            return this.data.size();
        endfunction // size   

        function automatic void make_random(int len, bit err=0);
            this.data = new [len];
            foreach ( this.data[i] ) begin
                this.data[i] = "a"+ $urandom() % ("z"-"a"+1);
            end
            this.err = err;
        endfunction // make_random      

 

        function automatic bit is_data_equal(ref data_t data_b );
            if (this.data.size() != data_b.size()) begin
                `LOG_ERROR( $sformatf("Packet data size mismatch match this.data.size=%0d, data_b.size=%0d.", this.data.size(), data_b.size()) );
                return 0;
            end 
            foreach ( this.data[i] ) begin
                if (this.data[i]!=data_b[i]) begin
                    `LOG_ERROR( $sformatf("Packet data mismatch this.data[%0d]=%0x, data_b[%0d]=%0x.",i, this.data[i], i, data_b[i]) );
                    return 0;
                end
            end
            return 1;
        endfunction // is_data_equal


        function automatic bit is_packet_equal(ref Packet pkt_b);

            if (this.err != pkt_b.err) begin
                `LOG_ERROR( $sformatf("Packet error mismatch this.err=%0b, pkt_b.err=%0b.",this.err, pkt_b.err) );
                return 0;
            end

            return this.is_data_equal(pkt_b.data);

        endfunction // is_packet_equal

    endclass



endpackage