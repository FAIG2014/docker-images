

package LCD_Controller_pkg;





endpackage
