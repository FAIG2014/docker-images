

package string_pkg;
	typedef byte string_t[16];



endpackage