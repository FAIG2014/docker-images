


module avalon_st_sink (input clk, interface.tx avalon_st);


endmodule