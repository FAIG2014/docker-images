module generic_top
    #( )
    (
        input               clk, 
        input               reset
    );


endmodule 
