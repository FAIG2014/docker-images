


module avalon_st_source (input clk, interface.tx avalon_st);


endmodule